 `define no_of_trans 20
 `define OP_WIDTH  8
 `define CMD_WIDTH  4

`define ROR_WIDTH                $clog2(`OP_WIDTH)

`define MAX ((1<<`OP_WIDTH)-1)
